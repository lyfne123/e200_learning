`include "e203_defines.v"

module e203_exu_alu_rglr(

);
endmodule